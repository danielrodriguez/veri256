
module padder1(in, byte_num, out);
    input      [543:0] in;
    input      [7:0]  byte_num;
    output reg [543:0] out;
    
    always @ (*)
      case (byte_num)
        0: out =               544'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        1: out = {in[543:536], 536'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        2: out = {in[543:528], 528'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        3: out = {in[543:520], 520'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        4: out = {in[543:512], 512'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        5: out = {in[543:504], 504'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        6: out = {in[543:496], 496'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        7: out = {in[543:488], 488'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        8: out = {in[543:480], 480'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        9: out = {in[543:472], 472'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        10: out = {in[543:464], 464'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        11: out = {in[543:456], 456'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        12: out = {in[543:448], 448'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        13: out = {in[543:440], 440'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        14: out = {in[543:432], 432'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        15: out = {in[543:424], 424'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        16: out = {in[543:416], 416'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        17: out = {in[543:408], 408'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        18: out = {in[543:400], 400'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        19: out = {in[543:392], 392'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        20: out = {in[543:384], 384'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        21: out = {in[543:376], 376'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        22: out = {in[543:368], 368'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        23: out = {in[543:360], 360'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        24: out = {in[543:352], 352'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        25: out = {in[543:344], 344'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        26: out = {in[543:336], 336'h010000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        27: out = {in[543:328], 328'h0100000000000000000000000000000000000000000000000000000000000000000000000000000000};
        28: out = {in[543:320], 320'h01000000000000000000000000000000000000000000000000000000000000000000000000000000};
        29: out = {in[543:312], 312'h010000000000000000000000000000000000000000000000000000000000000000000000000000};
        30: out = {in[543:304], 304'h0100000000000000000000000000000000000000000000000000000000000000000000000000};
        31: out = {in[543:296], 296'h01000000000000000000000000000000000000000000000000000000000000000000000000};
        32: out = {in[543:288], 288'h010000000000000000000000000000000000000000000000000000000000000000000000};
        33: out = {in[543:280], 280'h0100000000000000000000000000000000000000000000000000000000000000000000};
        34: out = {in[543:272], 272'h01000000000000000000000000000000000000000000000000000000000000000000};
        35: out = {in[543:264], 264'h010000000000000000000000000000000000000000000000000000000000000000};
        36: out = {in[543:256], 256'h0100000000000000000000000000000000000000000000000000000000000000};
        37: out = {in[543:248], 248'h01000000000000000000000000000000000000000000000000000000000000};
        38: out = {in[543:240], 240'h010000000000000000000000000000000000000000000000000000000000};
        39: out = {in[543:232], 232'h0100000000000000000000000000000000000000000000000000000000};
        40: out = {in[543:224], 224'h01000000000000000000000000000000000000000000000000000000};
        41: out = {in[543:216], 216'h010000000000000000000000000000000000000000000000000000};
        42: out = {in[543:208], 208'h0100000000000000000000000000000000000000000000000000};
        43: out = {in[543:200], 200'h01000000000000000000000000000000000000000000000000};
        44: out = {in[543:192], 192'h010000000000000000000000000000000000000000000000};
        45: out = {in[543:184], 184'h0100000000000000000000000000000000000000000000};
        46: out = {in[543:176], 176'h01000000000000000000000000000000000000000000};
        47: out = {in[543:168], 168'h010000000000000000000000000000000000000000};
        48: out = {in[543:160], 160'h0100000000000000000000000000000000000000};
        49: out = {in[543:152], 152'h01000000000000000000000000000000000000};
        50: out = {in[543:144], 144'h010000000000000000000000000000000000};
        51: out = {in[543:136], 136'h0100000000000000000000000000000000};
        52: out = {in[543:128], 128'h01000000000000000000000000000000};
        53: out = {in[543:120], 120'h010000000000000000000000000000};
        54: out = {in[543:112], 112'h0100000000000000000000000000};
        55: out = {in[543:104], 104'h01000000000000000000000000};
        56: out = {in[543:96], 96'h010000000000000000000000};
        57: out = {in[543:88], 88'h0100000000000000000000};
        58: out = {in[543:80], 80'h01000000000000000000};
        59: out = {in[543:72], 72'h010000000000000000};
        60: out = {in[543:64], 64'h0100000000000000};
        61: out = {in[543:56], 56'h01000000000000};
        62: out = {in[543:48], 48'h010000000000};
        63: out = {in[543:40], 40'h0100000000};
        64: out = {in[543:32], 32'h01000000};
        65: out = {in[543:24], 24'h010000};
        66: out = {in[543:16], 16'h0100};
        67: out = {in[543:8], 8'h01};
        default: out = 0;
      endcase
endmodule
