
module point_add_jaco_test;
reg clk, rst_n, start;
reg [255:0] px, py, pz, m;
reg [255:0] qx, qy, qz;
wire [255:0] rx, ry, rz;
wire ready;

    point_add_jaco inst (clk, rst_n, start, px, py, pz, qx, qy, qz, m, rx, ry, rz, ready);
    
    always #1 clk = ~ clk;

    initial begin
        clk = 0;
        rst_n = 0;
        start = 0;
    end

    initial begin

        #1;
        rst_n = 0;
        #5;
        rst_n = 1;
        m = 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f;
        px = 256'h6530e2c73e814654aca93bebcd0af877f23f209fec8751630869e6efed35e518;
        py = 256'hd5a7d0c22333b02db0a39e026e2d8bc08bfa96985b7385fcce36534283fd2a50;
        pz = 256'd68105346093711073138579907681248754787874622517682867538427217502358489265635;
        qx = 256'hfdbe15a370b1f0bfbab2c50f45fcffba4ddafe3fafc433471dd75b296592bb5d;
        qy = 256'hdce62b2b3d046deaa601ede644857dfc14e41e1f64418f62998b152c2092a61a;
        qz = 256'h60b3c4c75b3db9cabf9b9c03d327420bbb5bdb79b4ffd23d4f64a8f4f72f5f97;
        start = 1;
        #1
        while(!ready) 
          #1;
        // {'__name__': '__main__', '__doc__': None, '__package__': None, '__loader__': <_frozen_importlib_external.SourceFileLoader object at 0x1045a39e0>, '__spec__': None, '__annotations__': {}, '__builtins__': <module 'builtins' (built-in)>, '__file__': '/Users/drodriguez/src/veri/ecpt4o/ref_padd.py', '__cached__': None, 'random': <module 'random' from '/opt/homebrew/Cellar/python@3.12/3.12.3/Frameworks/Python.framework/Versions/3.12/lib/python3.12/random.py'>, 'm': 115792089237316195423570985008687907853269984665640564039457584007908834671663, 'verihex': <function verihex at 0x1045ace00>, 'mod': <function mod at 0x10462dc60>, 'double': <function double at 0x1046e8a40>, 'x1': 45769971532305571726516453356493850598853547143204083697208382823702101091608, 'y1': 96639141005230710270452256843679094305588790932055591848732050678161281460816, 'z1': 68105346093711073138579907681248754787874622517682867538427217502358489265635, 'x2': 114771000976887055740640413079191079519382180248934776414271382785218063809373, 'y2': 99915499454014124445154277383509266192157066822480400413009468884083769779738, 'z2': 43739657205511072834862987620297510373768801968260701592923611689706733920151, 'i1': 41354120465430223433051873631124625113762993905279795537365687481188842359957, 'i2': 58886910545427237629564241436743381634166202722033819623276003072070391878846, 'j1': 501601615292213631924076007461990473749032130170217725755094839061926825807, 'j2': 85670370135857526338133017495959951150852752677924580660025631604385419531169, 'u1': 63267789754937460876416011582716671501434725777759612516866937587665764096584, 'u2': 20220995530093652303813541378363213733674771260974530723171568937799392668296, 'h': 43046794224843808572602470204353457767759954516785081793695368649866371428288, 'f': 21429479383347542865612776619158301674632038561543049883444398670017659897753, 'k1': 79359341465883474679889964073936903534248609536557660965284185186566923060032, 'k2': 91172894517996927738770693539482592070104936587943853062644537276055647677264, 'v': 79487531048350101390060086977257843427623419988693181716388639095162082771770, 'g': 22711068145128009492520957964449068134531704953336680411036387437424560462836, 'r': 92164983133089289305809526077596530781557330562868179844736879828931385437199, 'x3': 72681894825567760862615927599087056320845441075635806264233766360389969293732, 'y3': 82809877791380838586607267121578203069865497243855582219939467962465479493853, 'z3': 25968162136531316409799580775230252462956021394676982819186909827493618081234, 'tmpx': 72778447635572795594131536226927469552311721741041618095876534896465493946, 'tmp2v': 43182972859384007356549188945827779001976855311745799393319694182415330871877, 'tmp2': 1969679410820158973543668274523428989131141230488957269204319490798067202147, 'tmp4': 34951890856755515810507386161633133772535628652273939088722435536241422379957, 'tmp5': 32139378633861144737346304156714511304920285935122190673527902310817799285157, 'tmp6': 100241031010857461062616115067868006747929196627313615160641690553259234238803, 'tmp7': 47690436860319879098301174097534412410261073973449139552343795765467399718017}
        check(256'ha0b07ea14e5e03b41a84a7532dd64f7ff2c8758f9ae69f94cc68612eeb10b1a4,
        256'hb714bad86a2585b2aad05781f5e1b55a17e6cf63e4384f8e1e60eb9a17cb08dd,
        256'h3969757b304ec0ed9652c0597be4def0042d5186f75db729cdceaf4c82855dd2);
        
        $display("✅ add 0x6530e2c73e814654aca93bebcd0af877f23f209fec8751630869e6efed35e518,0xdce62b2b3d046deaa601ede644857dfc14e41e1f64418f62998b152c2092a61a ok");
          
          

        #1;
        rst_n = 0;
        #5;
        rst_n = 1;
        m = 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f;
        px = 256'h8d6304e5ce442154f42d4eaac6094251aa16eb79be679933ec5c5534ffd1e92b;
        py = 256'h237c69a2387e0550d295256040016eece65bf1594b752b516f72291aef98aafb;
        pz = 256'd36123800115072815261167518527126549661538776391974639015416415736108496932162;
        qx = 256'h25df8eee371899cd6c7e9e32c42712e8825086942231de23747d2d0306ec4e24;
        qy = 256'h28129cc916f417cf429d4d3006cf7003bb231cbfe5ee1c79e940b3550f2cdc9e;
        qz = 256'h817f15fcc449bb207bd56c32c385bbfa11b9668eb0378cfe89269f58423c81b1;
        start = 1;
        #1
        while(!ready) 
          #1;
        // {'__name__': '__main__', '__doc__': None, '__package__': None, '__loader__': <_frozen_importlib_external.SourceFileLoader object at 0x1021c79e0>, '__spec__': None, '__annotations__': {}, '__builtins__': <module 'builtins' (built-in)>, '__file__': '/Users/drodriguez/src/veri/ecpt4o/ref_padd.py', '__cached__': None, 'random': <module 'random' from '/opt/homebrew/Cellar/python@3.12/3.12.3/Frameworks/Python.framework/Versions/3.12/lib/python3.12/random.py'>, 'm': 115792089237316195423570985008687907853269984665640564039457584007908834671663, 'verihex': <function verihex at 0x1021d0e00>, 'mod': <function mod at 0x102251c60>, 'double': <function double at 0x10230ca40>, 'x1': 63951063312189153972435565206907539583565780953660622426662867268014863149355, 'y1': 16050767793273946606552652819514558388038101199163562458174999733292429257467, 'z1': 36123800115072815261167518527126549661538776391974639015416415736108496932162, 'x2': 17130568763277283337321635906218481919661248549099711540580231559584322178596, 'y2': 18125399284293330333368214953310669934805337659208337719316035613233085471902, 'z2': 58572898795719601960342905452806406652454780246798982046433210768235171709361, 'i1': 62365985293682175807698104358492279207336930454934365212039320801695316281778, 'i2': 3252079316460830557507918159680856119303485286503071764817817120323078464677, 'j1': 4814025013790927517409240393469565733540015184311594232603443782143417986150, 'j2': 64678381036686259318952647541666240455026435454736325095741208138307007745042, 'u1': 80746565352782874356151423149546717253022537941887169337485318890123017324115, 'u2': 92955898044614661164530723396545218475366322287386390502682770965899211229392, 'h': 103582756545484408615191684761689406630926200320141342874260131932132640766386, 'f': 33203385803349891281385388306126823660650432189715140878324347911960209477846, 'k1': 100236567621809764729670687519570015343242073883597881616386903444564270808557, 'k2': 77548092568516084725982735321279019354207764253732344512442336150773962304752, 'v': 7869229424831306132920899131193457304928493683008435445148992523137262172819, 'g': 10976252762143921892483890896015782788775814158660234884632098106821498967475, 'r': 45376950106587360007375904396581991978068619259731074207889134587580617007610, 'x3': 5971453426651583065612438164842698943377923162928389924761003713428905231976, 'y3': 28669215681186805242413016724621941843321605536458924251443841141743763219454, 'z3': 69224248597147210654491052427881125349600115993068503295828127975871202377032, 'tmpx': 21709912276314195331454236427229613553234910528945260815058988759703429577614, 'tmp2v': 15738458849662612265841798262386914609856987366016870890297985046274524345638, 'tmp2': 110681997103747543705166890733386154944242669857883016723833510037000749437359, 'tmp4': 82012781422560738462753874008764213100921064321424092472389668895256986217905, 'tmp5': 60755719570375567799641508181388654215725957309379615825907156227140709009865, 'tmp6': 65618064610143006365206022518173135326640415741437436976857137922018394746455, 'tmp7': 110929744197548756858006470671903426742355526233582742888507602313031148935073}
        check(256'hd33b90dc96b6acc1203928ccfdd29aeecba6cf6b07fc2545d6058cd518f8668,
        256'h3f62337766822ac8ec2e8430a6f6190ac9ce8857439840f97280be29b7ae63fe,
        256'h990b8946bb876fd03804301f58c6c84a117e84eda60cf5573c59f9aa9fa6bd48);
        
        $display("✅ add 0x8d6304e5ce442154f42d4eaac6094251aa16eb79be679933ec5c5534ffd1e92b,0x28129cc916f417cf429d4d3006cf7003bb231cbfe5ee1c79e940b3550f2cdc9e ok");
          
          

        #1;
        rst_n = 0;
        #5;
        rst_n = 1;
        m = 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f;
        px = 256'h13d81646c12d69f8f54d0269dede060efaaeda5e8f5e85174019261245984689;
        py = 256'he5c461cfe7a553232d5fd51484db76ea6e84fc9894ffc29861bfa8fbf5ce93b9;
        pz = 256'd53619534275189359519343141123350208970985628933701644303988722354778453994320;
        qx = 256'h89f1ffc060fa2a2d73078303f93219a9bef8ee52e86a849b4e6eaf15181fb9d5;
        qy = 256'hd83eb405cc22ce3028a5b23ff0739c098fb2cf6c1ea233de49f27ab8f995cbf5;
        qz = 256'h7e8e8fc12bb8cbc997fdbff7363550ba4a735e091a1af4658bc30c5dfd0cd9;
        start = 1;
        #1
        while(!ready) 
          #1;
        // {'__name__': '__main__', '__doc__': None, '__package__': None, '__loader__': <_frozen_importlib_external.SourceFileLoader object at 0x1010ab9e0>, '__spec__': None, '__annotations__': {}, '__builtins__': <module 'builtins' (built-in)>, '__file__': '/Users/drodriguez/src/veri/ecpt4o/ref_padd.py', '__cached__': None, 'random': <module 'random' from '/opt/homebrew/Cellar/python@3.12/3.12.3/Frameworks/Python.framework/Versions/3.12/lib/python3.12/random.py'>, 'm': 115792089237316195423570985008687907853269984665640564039457584007908834671663, 'verihex': <function verihex at 0x1010b4e00>, 'mod': <function mod at 0x101135c60>, 'double': <function double at 0x1011f0a40>, 'x1': 8975736835034042996763297223645795222275875894427424260904915672329893725833, 'y1': 103926619424764315086054397476721009899496533853918081697675731056611220689849, 'z1': 53619534275189359519343141123350208970985628933701644303988722354778453994320, 'x2': 62394435530360169328965634633891917006907642162942632326635484529175203658197, 'y2': 97810362282641980974964684961381099050784798703915700947530510669183473535989, 'z2': 223606653758952509944401318355257933526266261903940143450097314200775625945, 'i1': 85667440800642460301481995318995168833601984448241598128417601377846631242979, 'i2': 95621977362891320765416300350955623911935196601744685036688306306974228569676, 'j1': 39366741035074937908286680201301304053492715534089567062139245288170001726302, 'j2': 33584790519998823683087766697001598419708389172150917959868534112808748833058, 'u1': 91227619196403472505959262359528761959816009340412958636249655619406557915421, 'u2': 54505550775472935424222193021127928294726177340771584033212276506476058639548, 'h': 36722068420930537081737069338400833665089831999641374603037379112930499275873, 'f': 64200167886680956097620644503930006082611369717434700544195825379212676014257, 'k1': 110667063161742393297373610262818526066060359286323380065122195016941778316980, 'k2': 58219477475201834846715977747739191121808505568856079036238103544981402013281, 'v': 100242800712335492385450487676734550298172030723642346858725736694164481059536, 'g': 86398207782746006461715324887112933998131124408078595156489638943811543789493, 'r': 104895171373081116901315265030158669888503707434934602057768182943920752607398, 'x3': 30149822837457663221670002261425865653991637496374442750639935662256095450159, 'y3': 97582186934429156035979797191782293673307606342322418109905403612500297959339, 'z3': 115685595423191064632989861330729898929245034562531830336802475543398365711579, 'tmpx': 114843335024812452568999992606207058397065714278018572428633825042676222897568, 'tmp2v': 84693512187354789347329990344781192743074076781644129677993889380420127447409, 'tmp2': 29994129619581546431505103550398536882367175557708056640071313921166280446901, 'tmp4': 48204031922468585819096291367304151062329553881026202569623494316574817159225, 'tmp5': 72670940038751585144027193145070803808425413020433434607053911595722889183102, 'tmp6': 65497328926217585643327310661262884892267196384345719125648323676912025140992, 'tmp7': 7173611112533999500699882483807918916158216636087715481405587918810864042110}
        check(256'h42a831eb1bbc3399063a6927b7f88872230fdd385f2abf5c849b586f49ab542f,
        256'hd7bd8f7fbf44cca20a387bb2a358363284f67047758deee6087be5b2f7cec7ab,
        256'hffc3ba04e57870a4c0f7cf9e71e9ce03c5bcdd931f88dd501bfc3fe3d626ccdb);
        
        $display("✅ add 0x13d81646c12d69f8f54d0269dede060efaaeda5e8f5e85174019261245984689,0xd83eb405cc22ce3028a5b23ff0739c098fb2cf6c1ea233de49f27ab8f995cbf5 ok");
          
          
        // mine, leave here
        #1;
        rst_n = 0;
        #10;
        rst_n = 1;
        m  = 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f;
        px = 256'hfed5b7e864ae24ed502e69af8acfe4c97190cbac30c2728c0d87afc60791219a;
        py = 256'h51898bfdf1b316664d1265ce8910b2177b522cdbf385e75f84c6059cdf3d0ca6;
        pz = 256'd1;
        qx = 256'hfd15b0a9c566cba7317e8c0826356ca9fd88cc6d49d48c180bded20418f92715;
        qy = 256'h7124f3c9f53b546921ab91834a6c099a6556abda6c89306c6ff86f48683a5645;
        qz = 256'ha31317fbe3662ccc9a24cb9d1221642ef6a459b7e70bcebf098c0b39be7a194c;
        start = 1;
        #1
        while(!ready) 
          #5;
        
        check(256'h660c64f81f03c2367e8bcaafb21c944cd28c2063065e4ac2c601d0fc7aa735fe,
        256'he7cbce74717c32a0a0d7c31d2666eada34078f59776d4e2cf7ac67221e412d34,
        256'h9f89ba13b552dd4fd47923330b225dfba18e6b0a48aca82c3052157763cf3176);

        $display("✅all good!");
        $finish;
    end

      task check;
        input [256:0] wishx, wishy, wishz;
        begin
          if (rx !== wishx)
            begin
              $display("❌ x actual: %0h", rx); 
              $display("❌ x expect: %0h", wishx); 
            end
          if (ry !== wishy)
            begin
              $display("❌ y actual: %0h ", ry);
              $display("❌ y expect: %0h", wishy); 
            end
          if (rz !== wishz)
            begin
              $display("❌ z actual: %0h", rz); 
              $display("❌ z expect: %0h", wishz); 
            end

            if (rx !== wishx | ry !== wishy | rz !== wishz)
              $finish;
        end
    endtask
endmodule
          
       
         
